module mod0(input i, output o);
endmodule