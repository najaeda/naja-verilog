`include "does_not_exist.v"

module should_not_parse ();
endmodule
