/*
  Unterminated pragma
*/

(* src = "/home/source/test.v"
module test();
endmodule