module mod0(input i0, output o0);
endmodule

module test(i, o, io);
  wire _i0_;
  wire _i1_;
  input i;
  wire i;
  output [3:0] o;
  wire [3:0] o;
  inout io;
  wire io;
endmodule