`include preprocess_include.v

module should_not_parse ();
endmodule
