module test10();

MOD
  // test:#
  // /home/foo/bar/elem.v:10
  // param0(1'b0)
  // param1('d0)
  // param2(1'b0)
  #(
   .elem10('d0)
  )
  ins (
   .INPUT1(1'b1)
  ,.INPUT2(1'b0)
  ,.INPUT3(1'b0)
  ,.INPUT4(1'b0)
);

endmodule