/*
  Focus on assign test
*/
module test(\asqrt[33] );
  wire n0, n1;

  assign n0 = n1;
  assign n1 = 1'b0;
endmodule