`include "preprocess_include_recursive.v"

module should_not_parse ();
endmodule
