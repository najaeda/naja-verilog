module test11();
//test octal

MOD
  #(
   .elem10('o0),
   .elem11(8'o84)
  )
  ins();

endmodule