` 
module empty_directive (input i, output o);
  wire w0;
  assign w0 = i;
  assign o = w0;
endmodule
