`include "include_unreadable.v"

module should_not_parse ();
endmodule
