`unknown_directive foo

module should_not_parse ();
endmodule
