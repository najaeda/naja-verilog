module test()
endmodule