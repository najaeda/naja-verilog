/*
  Syntax error
*/

module test();
  //Missing ";"
  model ins
endmodule