/*
  parameter assignments: string
*/
module test();
  mod #(
    .PARAM0(""),
    .PARAM1("A"),
    .PARAM2("VALUE")
  ) ins();
endmodule