`define

module should_not_parse ();
endmodule
