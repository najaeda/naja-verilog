/*
  Unterminated comment
*/

module test();
endmodule

/*
  This is not terminated