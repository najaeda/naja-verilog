`elsif SOME_FLAG

module should_not_parse ();
endmodule
