`include "unterminated_path

module should_not_parse ();
endmodule
