module mod1(input a, output b);
endmodule