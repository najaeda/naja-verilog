module test(input i);
endmodule
