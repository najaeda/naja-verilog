`timescale 1ns/1ps

module timescale_active (input i, output o);
  wire w0;
  assign w0 = i;
  assign o = w0;
endmodule
