`ifdef NEVER_CLOSED
module should_fail ();
endmodule
