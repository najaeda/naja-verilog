module test
endmodule
